//=============================================================================
// Release information
// Design version: sifive_sesame_rel3_190711
// Document version: OMC-V1.4-UG-R2.11, OMC-V1.4-IG-R1.00-SESAME
// Release generated at Thu Jul 11 15:30:19 2019
//=============================================================================

//=============================================================================
// Description :
// Generation time : 2019.06.27 on Thursday, 14:46:57
//=============================================================================


`ifndef __DOM_COG__CND_AXI_M0_DEFINE__
`define __DOM_COG__CND_AXI_M0_DEFINE__
  `define __ENABLE_AR_CH_RB_TOP_CHK__
  `define __ENABLE_AW_CH_RB_TOP_CHK__
  `define __ENABLE_R_CH_RB_TOP_CHK__
  `define __ENABLE_R_CH_RB_CORE_CHK__
`endif



// vim: tabstop=2 softtabstop=2 shiftwidth=2 expandtab autoindent smartindent
