//=============================================================================
// Release information
// Design version: sifive_sesame_rel3_190711
// Document version: OMC-V1.4-UG-R2.11, OMC-V1.4-IG-R1.00-SESAME
// Release generated at Thu Jul 11 15:30:19 2019
//=============================================================================

//=============================================================================
// Description :
// Generation time : 2019.06.27 on Thursday, 14:46:57
//=============================================================================


`ifndef __DOM_COG__SND_AXI_CTL_DEFINE__
`define __DOM_COG__SND_AXI_CTL_DEFINE__
  `define __ENABLE_DOM_COG__SND_AXI_CTL_CORE_CHK__
  `define __ENABLE_DOM_COG__SND_AXI_CTL_AR_TOP_CHK__
  `define __ENABLE_DOM_COG__SND_AXI_CTL_R_TOP_CHK__
  `define __ENABLE_DOM_COG__SND_AXI_CTL_AW_TOP_CHK__
  `define __ENABLE_DOM_COG__SND_AXI_CTL_W_TOP_CHK__
  `define __ENABLE_DOM_COG__SND_AXI_CTL_B_TOP_CHK__

`endif


// vim: tabstop=2 softtabstop=2 shiftwidth=2 expandtab autoindent smartindent
